module barrel_shifter
(
    input din[7:0],
    input shamt[2:0],
    input dir,
    input ari,

    output dout[7:0]
);





endmodule